module LED(
	input clk,
 

)



endmodule